`include "register.v"

//module random_access_memory #(parameter SIZE = 8)(input [SIZE-1:0] address, ) 
